.subckt TLine1
+a1 b1 c1 d1 e1 f1 ref1
+a2 b2 c2 d2 e2 f2 ref2

+length = 0.1016

.Model DEFAULT_2DEM_MODEL W MODELTYPE=RLGC N=6
+ L0=
+ 3.39704e-07
+ 2.50234e-08 3.38949e-07
+ 1.97042e-09 2.49640e-08 3.38945e-07
+ 1.55198e-10 1.96575e-09 2.49637e-08 3.38945e-07
+ 1.22242e-11 1.54832e-10 1.96575e-09 2.49640e-08 3.38949e-07
+ 9.65121e-13 1.22242e-11 1.55198e-10 1.97042e-09 2.50234e-08 3.39704e-07
+ C0=
+ 1.27267e-10
+ -9.33008e-12 1.28229e-10
+ -3.98550e-14 -9.32574e-12 1.28229e-10
+ -0.00000e+00 -4.04054e-14 -9.32574e-12 1.28229e-10
+ -0.00000e+00 -0.00000e+00 -4.04054e-14 -9.32574e-12 1.28229e-10
+ -0.00000e+00 -0.00000e+00 -0.00000e+00 -3.98550e-14 -9.33008e-12 1.27267e-10
+ R0=
+ 1.08362e+01
+ 0.00000e+00 1.08362e+01
+ 0.00000e+00 0.00000e+00 1.08362e+01
+ 0.00000e+00 0.00000e+00 0.00000e+00 1.08362e+01
+ 0.00000e+00 0.00000e+00 0.00000e+00 0.00000e+00 1.08362e+01
+ 0.00000e+00 0.00000e+00 0.00000e+00 0.00000e+00 0.00000e+00 1.08362e+01
+ G0=
+ 0.00000e+00
+ 0.00000e+00 0.00000e+00
+ 0.00000e+00 0.00000e+00 0.00000e+00
+ 0.00000e+00 0.00000e+00 0.00000e+00 0.00000e+00
+ 0.00000e+00 0.00000e+00 0.00000e+00 0.00000e+00 0.00000e+00
+ 0.00000e+00 0.00000e+00 0.00000e+00 0.00000e+00 0.00000e+00 0.00000e+00
+ Rs=
+ 1.62251e-03
+ 0.00000e+00 1.62251e-03
+ 0.00000e+00 0.00000e+00 1.62251e-03
+ 0.00000e+00 0.00000e+00 0.00000e+00 1.62251e-03
+ 0.00000e+00 0.00000e+00 0.00000e+00 0.00000e+00 1.62251e-03
+ 0.00000e+00 0.00000e+00 0.00000e+00 0.00000e+00 0.00000e+00 1.62251e-03
+ Gd=
+ 1.81717e-11
+ -1.26029e-12 1.82943e-11
+ 0.00000e+00 -1.26029e-12 1.82943e-11
+ 0.00000e+00 0.00000e+00 -1.26029e-12 1.82943e-11
+ 0.00000e+00 0.00000e+00 0.00000e+00 -1.26029e-12 1.82943e-11
+ 0.00000e+00 0.00000e+00 0.00000e+00 0.00000e+00 -1.26029e-12 1.81717e-11

W1 a1 b1 c1 d1 e1 f1 ref1 a2 b2 c2 d2 e2 f2 ref2
+ N=6 L='length' RLGCModel=DEFAULT_2DEM_MODEL FGD=0.00000e+00
.ENDS
