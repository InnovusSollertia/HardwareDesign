.subckt VRM pwr ngnd

+ Voltage = 0.9          $ Nominal Voltage

* power supply
Vsupply pwr ngnd 'Voltage'

.ends VRM
