

.subckt TL2 1 3 2 4 ngnd


WTL1 1 3 ngnd 2 4 ngnd n=2 RLGCfile=MTL_Z50000_ZD100000_V14224_VD14224_7.rlc
+ l=0.07112




.ends TL2
